module WorkingRam
(
   input clk, ce2Hd,
   input [15:0] BA,
   input SRAMn, BRWn,
   //input [8:0] hcount,
   //input BUF1BUF2n,
   
   input [7:0] data_to_sram,
   output [7:0] data_from_sram  
);
   
wire [10:0] addr = BA[11:1];        // TODO multiplex with hcount

wire WE6B = ~SRAMn & BA[0] & ~BRWn & ce2Hd;
wire WE6D = ~SRAMn & ~BA[0] & ~BRWn & ce2Hd;

wire [7:0] data_from_6B, data_from_6D;

sram #(.INIT_FILE("empty2k.ram")) ic6B
(
   .clk(clk),
   .we(WE6B),
   .addr(addr), 
   .din(data_to_sram),
   .dout(data_from_6B)
);

sram #(.INIT_FILE("empty2k.ram")) ic6D
(
   .clk(clk),
   .we(WE6D),
   .addr(addr), 
   .din(data_to_sram),
   .dout(data_from_6D)
);

assign data_from_sram = BA[0] ? data_from_6B : data_from_6D;

endmodule

